module get_target_number(input logic [2:0] counter, output logic [3:0] target_digit_1, target_digit_2, target_digit_3);



endmodule